`include "settings.h"

module Conditin_Check
(
    input  [3:0] condition,
    input  [3:0] status_register,
    output       condition_state
);

endmodule